`timescale 1ns/1ns

module XOR2_1bit(A, B, Out);

input A, B;
output Out;

assign #5 Out = A ^ B;

endmodule

module TB_XOR2_1bit();

reg A, B;
wire Out;

XOR2_1bit XOR(.A(A), .B(B), .Out(Out));

initial begin
	A = 1'b0; B = 1'b0;
	#100;
	A = 1'b0; B = 1'b1;
	#100;
	A = 1'b1; B = 1'b0;
	#100;
	A = 1'b1; B = 1'b1;
end
endmodule
