`timescale 1ns/1ns

module Mux64to1_4bit(I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, I32,
		     I33, I34, I35, I36, I37, I38, I39, I40, I41, I42, I43, I44, I45, I46, I47, I48, I49, I50, I51, I52, I53, I54, I55, I56, I57, I58, I59, I60, I61, I62, I63, Sel, Out);

input [3:0] I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, I32, I33, 
	    I34, I35, I36, I37, I38, I39, I40, I41, I42, I43, I44, I45, I46, I47, I48, I49, I50, I51, I52, I53, I54, I55, I56, I57, I58, I59, I60, I61, I62, I63;
input [5:0] Sel;
output [3:0] Out;

wire [3:0] tmp0, tmp1;

Mux32to1_4bit MUX0(.I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .I5(I5), .I6(I6), .I7(I7), .I8(I8), .I9(I9), .I10(I10), .I11(I11), .I12(I12), .I13(I13), .I14(I14),
		   .I15(I15), .I16(I16), .I17(I17), .I18(I18), .I19(I19), .I20(I20), .I21(I21), .I22(I22), .I23(I23), .I24(I24), .I25(I25), .I26(I26), .I27(I27),
		   .I28(I28), .I29(I29), .I30(I30), .I31(I31), .Sel(Sel[4:0]), .Out(tmp0));
Mux32to1_4bit MUX1(.I0(I32), .I1(I33), .I2(I34), .I3(I35), .I4(I36), .I5(I37), .I6(I38), .I7(I39), .I8(I40), .I9(I41), .I10(I42), .I11(I43), .I12(I44), .I13(I45), 
		   .I14(I46), .I15(I47), .I16(I48), .I17(I49), .I18(I50), .I19(I51), .I20(I52), .I21(I53), .I22(I54), .I23(I55), .I24(I56), .I25(I57), .I26(I58), 
		   .I27(I59), .I28(I60), .I29(I61), .I30(I62), .I31(I63), .Sel(Sel[4:0]), .Out(tmp1));

Mux2to1_4bit MUXOUT(.I0(tmp0), .I1(tmp1), .Sel(Sel[5]), .Out(Out));

endmodule
