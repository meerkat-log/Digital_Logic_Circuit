`timescale 1ns/1ns

module Comparator_32bit(A, B, ALB, AEB, AGB);

input [31:0] A, B;
output ALB, AEB, AGB;

wire CMP0_ALB, CMP1_ALB, CMP2_ALB, CMP3_ALB, CMP4_ALB, CMP5_ALB, CMP6_ALB;
wire CMP0_AEB, CMP1_AEB, CMP2_AEB, CMP3_AEB, CMP4_AEB, CMP5_AEB, CMP6_AEB;
wire CMP0_AGB, CMP1_AGB, CMP2_AGB, CMP3_AGB, CMP4_AGB, CMP5_AGB, CMP6_AGB;

Comparator_4bit CMP0(.A(A[3:0]), .B(B[3:0]), .ALBI(1'b0), .AEBI(1'b1), .AGBI(1'b0), .ALBO(CMP0_ALB), .AEBO(CMP0_AEB), .AGBO(CMP0_AGB));
Comparator_4bit CMP1(.A(A[7:4]), .B(B[7:4]), .ALBI(CMP0_ALB), .AEBI(CMP0_AEB), .AGBI(CMP0_AGB), .ALBO(CMP1_ALB), .AEBO(CMP1_AEB), .AGBO(CMP1_AGB));
Comparator_4bit CMP2(.A(A[11:8]), .B(B[11:8]), .ALBI(CMP1_ALB), .AEBI(CMP1_AEB), .AGBI(CMP1_AGB), .ALBO(CMP2_ALB), .AEBO(CMP2_AEB), .AGBO(CMP2_AGB));
Comparator_4bit CMP3(.A(A[15:12]), .B(B[15:12]), .ALBI(CMP2_ALB), .AEBI(CMP2_AEB), .AGBI(CMP2_AGB), .ALBO(CMP3_ALB), .AEBO(CMP3_AEB), .AGBO(CMP3_AGB));
Comparator_4bit CMP4(.A(A[19:16]), .B(B[19:16]), .ALBI(CMP3_ALB), .AEBI(CMP3_AEB), .AGBI(CMP3_AGB), .ALBO(CMP4_ALB), .AEBO(CMP4_AEB), .AGBO(CMP4_AGB));
Comparator_4bit CMP5(.A(A[23:20]), .B(B[23:20]), .ALBI(CMP4_ALB), .AEBI(CMP4_AEB), .AGBI(CMP4_AGB), .ALBO(CMP5_ALB), .AEBO(CMP5_AEB), .AGBO(CMP5_AGB));
Comparator_4bit CMP6(.A(A[27:24]), .B(B[27:24]), .ALBI(CMP5_ALB), .AEBI(CMP5_AEB), .AGBI(CMP5_AGB), .ALBO(CMP6_ALB), .AEBO(CMP6_AEB), .AGBO(CMP6_AGB));
Comparator_4bit CMP7(.A(A[31:28]), .B(B[31:28]), .ALBI(CMP6_ALB), .AEBI(CMP6_AEB), .AGBI(CMP6_AGB), .ALBO(ALB), .AEBO(AEB), .AGBO(AGB));

endmodule

module TB_Comparator_32bit();

reg [31:0] A, B;
wire ALB, AEB, AGB;

Comparator_32bit CMP(.A(A), .B(B), .ALB(ALB), .AEB(AEB), .AGB(AGB));

initial begin
	A = 32'H00000000; B = 32'H00000000;
	#300;
	A = 32'H00000000; B = 32'H00000001;
	#300;
	A = 32'H00000001; B = 32'H00000000;
	#300;
	A = 32'H00000001; B = 32'H00000001;
end
endmodule

